/*
 * SPI interface for MIPSfpga
 */

module mfp_ahb_spi(
           input        clk,
           input        resetn,
           input [7:0]  data,
           input        send,
           output       done,
           output       sdo,
           output       sck);

  // Add code here.

endmodule

 
