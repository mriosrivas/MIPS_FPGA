/*
 * Buzzer hardware for MIPSfpga
 */

module mipsfpga_ahb_buzzer(
              input        clk,
              input        resetn,
              input [31:0] numMicros,
              output       buzz);

  // Add code here.

endmodule

 
