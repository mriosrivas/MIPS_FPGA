// 
// mfp_config.vh
//
// Configuration settings for MIPSfpga
// 

`define MFP_USE_SLOW_CLOCK
`define MFP_INTERRUPTS
`define MFP_DEMO_CACHE_HITS_MISSES