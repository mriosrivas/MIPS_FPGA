/*
 * Seven-segment display timer for the Nexys4 DDR board
 *
 * January 25, 2017
 */

module mfp_ahb_sevensegtimer(
                     input            clk,
                     input            resetn,
                     input     [ 7:0] EN,
                     input     [31:0] DIGITS,
                     output    [ 7:0] DISPENOUT,
                     output    [ 6:0] DISPOUT);

    // add code here.
	
endmodule


