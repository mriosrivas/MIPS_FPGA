/*
 * Seven-segment display decoder
 *
 * January 25, 2017
 */

module mfp_ahb_sevensegdec(input      [3:0] data,
                           output reg [6:0] seg);

    // add code here.
	
endmodule
